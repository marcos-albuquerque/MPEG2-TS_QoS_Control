module mux_sync (
    input  wire [3:0]  sync,
    input  wire [1:0]  mux_ctrl,
    input  wire        en_mux,
    output reg         sync_out
);
    always @(*) begin
        if (en_mux) begin
            case (mux_ctrl)
                2'b00: sync_out = sync[0];
                2'b01: sync_out = sync[1];
                2'b10: sync_out = sync[2];
                2'b11: sync_out = sync[3];
                default: sync_out = 1'b0;
            endcase
        end else begin
            sync_out = 1'b0;
        end
    end
endmodule